// ZICBOM Cache-block management instructions.
//CBO_CLEAN,
//CBO_FLUSH,
//CBO_INVAL,
`DEFINE_INSTR(CBO_CLEAN,   I_FORMAT, SYSTEM, RV64ZICBOM)
`DEFINE_INSTR(CBO_FLUSH,   I_FORMAT, SYSTEM, RV64ZICBOM)
`DEFINE_INSTR(CBO_INVAL,   I_FORMAT, SYSTEM, RV64ZICBOM)

