// Already implemented -ZVKT Vector data-independent execution latency
//VCLMUL_VV ,
//VCLMUL_VX ,
//VCLMULH_VV,
//VCLMULH_VX,

