// ZIMOP may-be-operations
//MOP_R_N   , 
//MOP_RR_N  ,

`DEFINE_INSTR(MOP_R_N  ,   R_FORMAT, SYSTEM, RV64ZIMOP)
`DEFINE_INSTR(MOP_RR_N  ,   R_FORMAT, SYSTEM, RV64ZIMOP)

