// ZICBOP Cache-block prefetch instructions
//PREFETCH_I,
//PREFETCH_R,
//PREFETCH_W,
`DEFINE_INSTR(PREFETCH_I,   I_FORMAT, SYSTEM, RV64ZICBOP)
`DEFINE_INSTR(PREFETCH_R,   I_FORMAT, SYSTEM, RV64ZICBOP)
`DEFINE_INSTR(PREFETCH_W,   I_FORMAT, SYSTEM, RV64ZICBOP)

