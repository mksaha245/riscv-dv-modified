// ZVBB  Vector basic bit-manipulation instructionS
    //VANDN_VV , 
    //VANDN_VX , 
    //VBREV_V  ,
    //VBREV8_V ,
    //VREV8_V  ,
    //VCLZ_V   ,
    //VCTZ_V   ,
    //VCOPOP_V , 
    //VROL_VV  ,
    //VROL_VX  ,
    //VROR_VV  ,
    //VROR_VX  ,
    //VROR_VI  ,
    //VWSLL_VV , 
    //VWSLL_VX , 
    //VWSLL_VI , 

`DEFINE_VA_INSTR(VANDN_VV,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VANDN_VX,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VBREV_V  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VBREV8_V ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VREV8_V  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VCLZ_V   ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VCTZ_V   ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VCOPOP_V ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VROL_VV  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VROL_VX  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VROR_VV  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VROR_VX  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VROR_VI  ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX},UIMM)
`DEFINE_VA_INSTR(VWSLL_VV ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VWSLL_VX ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX})
`DEFINE_VA_INSTR(VWSLL_VI ,     VA_FORMAT, ARITHMETIC, RV64ZVBB, {VV, VX},UIMM)

