`DEFINE_B_INSTR(SM4ED,  	R_FORMAT, ARITHMETIC, RV64ZKSED, UIMM)
`DEFINE_B_INSTR(SM4KS,  	R_FORMAT, ARITHMETIC, RV64ZKSED, UIMM)

