// ZAWRS Wait-on-reservation-set instructions
//WRS_NTO    ,
//WRS_STO    ,
`DEFINE_INSTR(WRS_NTO,   I_FORMAT, SYSTEM, RV64ZIHINTPAUSE)
`DEFINE_INSTR(WRS_STO,   I_FORMAT, SYSTEM, RV64ZIHINTPAUSE)

