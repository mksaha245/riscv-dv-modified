// ZICOND Integer conditional operations
//CZERO_EQZ
//CZERO_NEZ

`DEFINE_INSTR(CZERO_EQZ  ,   R_FORMAT, ARITHMETIC, RV64ZICOND)
`DEFINE_INSTR(CZERO_NEZ  ,   R_FORMAT, ARITHMETIC, RV64ZICOND)

