/*/ ZCB Additional compressed instructions
    C_LBU     ,  
    C_LHU     ,
    C_LH      ,
    C_SB      ,
    C_SH      ,
    C_ZEXT_B  ,
    C_SEXT_B  ,
    C_ZEXT_H  ,
    C_SEXT_H  ,
    C_ZEXT_W  ,
    C_NOT     ,
    C_MUL     ,
*/

`DEFINE_INSTR(C_LBU      ,   CL_FORMAT, LOAD, RV64ZCB)
`DEFINE_INSTR(C_LHU      ,   CL_FORMAT, LOAD, RV64ZCB)
`DEFINE_INSTR(C_LH       ,   CL_FORMAT, LOAD, RV64ZCB)
`DEFINE_INSTR(C_SB       ,   CS_FORMAT, STORE, RV64ZCB)
`DEFINE_INSTR(C_SH       ,   CS_FORMAT, STORE, RV64ZCB)
`DEFINE_INSTR(C_ZEXT_B   ,   CR_FORMAT, ARITHMETIC, RV64ZCB)
`DEFINE_INSTR(C_SEXT_B   ,   CR_FORMAT, ARITHMETIC, RV64ZCB)
`DEFINE_INSTR(C_ZEXT_H   ,   CR_FORMAT, ARITHMETIC, RV64ZCB)
`DEFINE_INSTR(C_SEXT_H   ,   CR_FORMAT, ARITHMETIC, RV64ZCB)
`DEFINE_INSTR(C_ZEXT_W   ,   CR_FORMAT, ARITHMETIC, RV64ZCB)
`DEFINE_INSTR(C_NOT      ,   CR_FORMAT, ARITHMETIC, RV64ZCB)
`DEFINE_INSTR(C_MUL      ,   CR_FORMAT, ARITHMETIC, RV64ZCB)

