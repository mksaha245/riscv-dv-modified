/*
 * Modified by Mukesh
 * Adding instruction for RV16FH exntension
 * Floating Point Half Prescision
 *
 */

`DEFINE_FP_INSTR(FLH      ,I_FORMAT, LOAD, RV16FH)
`DEFINE_FP_INSTR(FSH      ,S_FORMAT, STORE, RV16FH)
`DEFINE_FP_INSTR(FMADD_H  ,R4_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FMSUB_H  ,R4_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FNMSUB_H ,R4_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FNMADD_H ,R4_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FADD_H   ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FSUB_H   ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FMUL_H   ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FDIV_H   ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FSQRT_H  ,I_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FSGNJ_H  ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FSGNJN_H ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FSGNJX_H ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FMIN_H   ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FMAX_H   ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FEQ_H    ,R_FORMAT, COMPARE, RV16FH)
`DEFINE_FP_INSTR(FLT_H    ,R_FORMAT, COMPARE, RV16FH)
`DEFINE_FP_INSTR(FLE_H    ,R_FORMAT, COMPARE, RV16FH)
`DEFINE_FP_INSTR(FCLASS_H ,R_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FMV_X_H  ,I_FORMAT, ARITHMETIC, RV16FH)
`DEFINE_FP_INSTR(FMV_H_X  ,I_FORMAT, ARITHMETIC, RV16FH)

