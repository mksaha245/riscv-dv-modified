`DEFINE_B_INSTR(SHA256SIG0, R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA256SIG1, R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA256SUM0, R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA256SUM1, R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA512SIG0,R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA512SIG1,R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA512SUM0,R_FORMAT, ARITHMETIC, RV64ZKNH)
`DEFINE_B_INSTR(SHA512SUM1,R_FORMAT, ARITHMETIC, RV64ZKNH)

