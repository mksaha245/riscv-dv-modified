// ZVFHMIN Vector Minimal Half-precision floating-point
//VFNCVT_F_F_V,
//VFWCVT_F_F_W,
