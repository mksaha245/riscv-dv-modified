/*/ ZCMOP  Compressed may-be-operations
    C_MOP_1   , 
    C_MOP_3   ,
    C_MOP_5   ,
    C_MOP_7   ,
    C_MOP_9   ,
    C_MOP_11  ,
    C_MOP_13  ,
    C_MOP_15  ,
*/

`DEFINE_INSTR(C_MOP_1   ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_3   ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_5   ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_7   ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_9   ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_11  ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_13  ,   R_FORMAT, SYSTEM, RV64ZCMOP)
`DEFINE_INSTR(C_MOP_15  ,   R_FORMAT, SYSTEM, RV64ZCMOP)

