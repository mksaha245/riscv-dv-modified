`DEFINE_B_INSTR(AES64DS,  R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(AES64DSM, R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(AES64IM,  R_FORMAT, ARITHMETIC, RV64ZBK)

`DEFINE_B_INSTR(AES64ES,  R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(AES64ESM, R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(AES64KS1I,I_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(AES64KS2, R_FORMAT, ARITHMETIC, RV64ZBK)

`DEFINE_B_INSTR(SHA256SIG0, R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA256SIG1, R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA256SUM0, R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA256SUM1, R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA512SIG0,R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA512SIG1,R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA512SUM0,R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SHA512SUM1,R_FORMAT, ARITHMETIC, RV64ZBK)

`DEFINE_B_INSTR(SM4ED,  	R_FORMAT, ARITHMETIC, RV64ZBK, UIMM)
`DEFINE_B_INSTR(SM4KS,  	R_FORMAT, ARITHMETIC, RV64ZBK, UIMM)

`DEFINE_B_INSTR(SM3P0,  	R_FORMAT, ARITHMETIC, RV64ZBK)
`DEFINE_B_INSTR(SM3P1,  	R_FORMAT, ARITHMETIC, RV64ZBK)

//`DEFINE_B_INSTR(SHA512SIG0H,R_FORMAT, ARITHMETIC, RV64ZBK)
//`DEFINE_B_INSTR(SHA512SIG0L,R_FORMAT, ARITHMETIC, RV64ZBK)
//`DEFINE_B_INSTR(SHA512SIG1H,R_FORMAT, ARITHMETIC, RV64ZBK)
//`DEFINE_B_INSTR(SHA512SIG1L,R_FORMAT, ARITHMETIC, RV64ZBK)
//`DEFINE_B_INSTR(SHA512SUM0R,R_FORMAT, ARITHMETIC, RV64ZBK)
//`DEFINE_B_INSTR(SHA512SUM1R,R_FORMAT, ARITHMETIC, RV64ZBK)

