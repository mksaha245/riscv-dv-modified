`DEFINE_B_INSTR(SM3P0,  	R_FORMAT, ARITHMETIC, RV64ZKSH)
`DEFINE_B_INSTR(SM3P1,  	R_FORMAT, ARITHMETIC, RV64ZKSH)

