// ZIHINTNTL Non-temporal locality hints.
//NTL_P1    , 
//NTL_PALL  ,
//NTL_S1    ,
//NTL_ALL   ,

`DEFINE_INSTR(NTL_P1  ,   I_FORMAT, ARITHMETIC, RV64ZIHINTPAUSE)
`DEFINE_INSTR(NTL_PALL,   I_FORMAT, ARITHMETIC, RV64ZIHINTPAUSE)
`DEFINE_INSTR(NTL_S1  ,   I_FORMAT, ARITHMETIC, RV64ZIHINTPAUSE)
`DEFINE_INSTR(NTL_ALL ,   I_FORMAT, ARITHMETIC, RV64ZIHINTPAUSE)

