/*
 * Copyright 2018 Google LLC
 * Copyright 2021 Silicon Labs, Inc.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`DEFINE_B_INSTR(CLMUL,  R_FORMAT, ARITHMETIC, RV64ZBKC)
`DEFINE_B_INSTR(CLMULH,  R_FORMAT, ARITHMETIC, RV64ZBKC)
`DEFINE_B_INSTR(CLMULR,  R_FORMAT, ARITHMETIC, RV64ZBKC)

`DEFINE_B_INSTR(CLMUL_W,  R_FORMAT, ARITHMETIC, RV64ZBKC)
`DEFINE_B_INSTR(CLMULH_W, R_FORMAT, ARITHMETIC, RV64ZBKC)
`DEFINE_B_INSTR(CLMULR_W, R_FORMAT, ARITHMETIC, RV64ZBKC)

